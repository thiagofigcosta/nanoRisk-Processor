module nRProcessor(clk,reset);

  input clk,reset;
  wire[7:0] im_addr,im_out;
  wire[7:0] dm_out;
  wire[7:0] nxtmux_in0,nxtmux_in1;
  wire[7:0] ctrlmux1_in0;
  wire nxtmux_sel,ctrlmux2_sel;
  wire ctrl2Cmp_out;
  wire adder_input;
  wire ULA_Zer0,branchAND_out;
  wire[1:0] regs_ovrflw;
  wire[7:0] regs_in0;
  wire[3:0] regs_adrIn0,regs_adrOut1;
  wire[7:0] regs_out0,regs_out1,regs_out2;
  wire[7:0] nxt_in;
  wire[7:0] ghost0_in,ghost1_in,ghost0_out,ghost1_out;
  wire ctrl_tmpwr,ctrl_hlt,ctrl_jmp,ctrl_brc,ctrl_rgr,ctrl_ala;
  wire[1:0] ctrl_rgw;
  wire[3:0] ctrl_alo,ctrl_ioc;
  wire[7:0] ULA_in1,ULA_out;
  wire haltNOTscape,haltScape;
  wire realClk,bitshift_out0;
  
  
  nR_Memory InstructionsMemory(clk,8'b00000000,im_out,8'b00000000,im_addr,1'b0,1'b1,1'b0); 
  nR_Register Next(clk,nxt_in,im_addr,reset);
  nR_Memory DataMemory(realClk,regs_out1,dm_out,ULA_out,ULA_out,ctrl_ioc[1],ctrl_ioc[0],1'b0); 
  nR_MUX2 NextMUX(nxtmux_in0,nxtmux_in1,nxtmux_sel,nxt_in);
  nR_FluxCtrl FluxControl(branchAND_out,ctrl_jmp,nxtmux_sel);
  nR_AND2 FluxAND(ctrl_brc,ULA_Zer0,branchAND_out);
  nR_OR4 AdderOr(reset,ctrl_hlt,haltScape,1'b0,adder_input);
  nR_Adder Adder(im_addr,{7'b0,adder_input},nxtmux_in0);
  nR_BitShifter BitShift(clk,bitshift_out0,realClk,1'b0);
  nR_8AND2 Ghost0_And(im_out,bitshift_out0,ghost0_in);
  nR_8AND2 Ghost1_And(im_out,realClk,ghost1_in);
  nR_Register Ghost0(clk,ghost0_in,ghost0_out,reset);
  nR_Register Ghost1(clk,ghost1_in,ghost1_out,reset);
  nR_MUX2 CtrlMUX1(ctrlmux1_in0,regs_out2,ctrl_brc,nxtmux_in1);
  nR_MUX2 CtrlMUX2(ghost1_out,regs_out1,ctrlmux2_sel,ctrlmux1_in0);
  nR_BitCmp Ctrl2Cmp(ghost1_out,ctrl2Cmp_out);
  nR_NOT Ctrl2Not(ctrl2Cmp_out,ctrlmux2_sel);
  nR_Control Control(realClk,ghost0_out[7:4],ctrl_tmpwr,ctrl_hlt,ctrl_jmp,ctrl_brc,ctrl_rgw,ctrl_ioc,ctrl_rgr,ctrl_alo,ctrl_ala);
  nR_MUX2 RegWriteMUX(8'b00000010,{4'b0,ghost0_out[3:0]},ctrl_tmpwr,regs_adrIn0);
  nR_RegisterBank Registers(realClk,regs_in0,regs_out0,regs_out1,regs_out2,regs_adrIn0,ghost1_out[7:4],regs_adrOut1,ghost1_out[3:0],ctrl_ioc[3],ctrl_ioc[2],reset,regs_ovrflw);
  nR_MUX2 AdrRead1MUX({4'b0,ghost0_out[3:0]},{4'b0,ghost1_out[3:0]},ctrl_rgr,regs_adrOut1);
  nR_MUX4 WriteMUX(ULA_out,nxtmux_in0,dm_out,ghost1_out,ctrl_rgw,regs_in0);
  nR_MUX2 ALUMUX(regs_out1,{4'b0,ghost1_out[3:0]},ctrl_ala,ULA_in1);
  nR_ALU ULALA(regs_out0,ULA_in1,ctrl_alo,ULA_Zer0,ULA_out,regs_ovrflw);
  nR_BitCmp HaltCmp(regs_out1,haltNOTscape);
  nR_NOT HaltNot(haltNOTscape,haltScape);
  
  always@(reset) begin 
    DataMemory.m_mem[0]<=8'b00000001;
	DataMemory.m_mem[1]<=8'b00101100;
	DataMemory.m_mem[2]<=8'b00000000;
	DataMemory.m_mem[3]<=8'b10010110;
	DataMemory.m_mem[4]<=8'b00000010;
	DataMemory.m_mem[5]<=8'b10011010;
	DataMemory.m_mem[6]<=8'b00000001;
	DataMemory.m_mem[7]<=8'b01100101;
	DataMemory.m_mem[8]<=8'b00000000;
	DataMemory.m_mem[9]<=8'b11011100;
	DataMemory.m_mem[10]<=8'b00000001;
	DataMemory.m_mem[11]<=8'b11100000;
	DataMemory.m_mem[12]<=8'b00000001;
	DataMemory.m_mem[13]<=8'b00010100;
	DataMemory.m_mem[14]<=8'b00000010;
	DataMemory.m_mem[15]<=8'b10011010;
	DataMemory.m_mem[16]<=8'b00000001;
	DataMemory.m_mem[17]<=8'b00000001;
	DataMemory.m_mem[18]<=8'b00000010;
	DataMemory.m_mem[19]<=8'b00000010;
	DataMemory.m_mem[20]<=8'b00001000;
	DataMemory.m_mem[21]<=8'b00101000;
	DataMemory.m_mem[22]<=8'b00011010;
	DataMemory.m_mem[23]<=8'b00011100;
	DataMemory.m_mem[24]<=8'b00010000;
  end
  
initial begin
#1 begin
//data seg
	DataMemory.m_mem[0]<=8'b00000001;
	DataMemory.m_mem[1]<=8'b00101100;
	DataMemory.m_mem[2]<=8'b00000000;
	DataMemory.m_mem[3]<=8'b10010110;
	DataMemory.m_mem[4]<=8'b00000010;
	DataMemory.m_mem[5]<=8'b10011010;
	DataMemory.m_mem[6]<=8'b00000001;
	DataMemory.m_mem[7]<=8'b01100101;
	DataMemory.m_mem[8]<=8'b00000000;
	DataMemory.m_mem[9]<=8'b11011100;
	DataMemory.m_mem[10]<=8'b00000001;
	DataMemory.m_mem[11]<=8'b11100000;
	DataMemory.m_mem[12]<=8'b00000001;
	DataMemory.m_mem[13]<=8'b00010100;
	DataMemory.m_mem[14]<=8'b00000010;
	DataMemory.m_mem[15]<=8'b10011010;
	DataMemory.m_mem[16]<=8'b00000001;
	DataMemory.m_mem[17]<=8'b00000001;
	DataMemory.m_mem[18]<=8'b00000010;
	DataMemory.m_mem[19]<=8'b00000010;
	DataMemory.m_mem[20]<=8'b00001000;
	DataMemory.m_mem[21]<=8'b00101000;
	DataMemory.m_mem[22]<=8'b00011010;
	DataMemory.m_mem[23]<=8'b00011100;
	DataMemory.m_mem[24]<=8'b00010000;

//instructions seg
	InstructionsMemory.m_mem[0]<=8'b11000111;
	InstructionsMemory.m_mem[1]<=8'b00010001;
	InstructionsMemory.m_mem[2]<=8'b11001000;
	InstructionsMemory.m_mem[3]<=8'b00010101;
	InstructionsMemory.m_mem[4]<=8'b11100111;
	InstructionsMemory.m_mem[5]<=8'b00000111;
	InstructionsMemory.m_mem[6]<=8'b11101000;
	InstructionsMemory.m_mem[7]<=8'b00001000;
	InstructionsMemory.m_mem[8]<=8'b11010010;
	InstructionsMemory.m_mem[9]<=8'b10001010;
	InstructionsMemory.m_mem[10]<=8'b10110010;
	InstructionsMemory.m_mem[11]<=8'b00000000;
	InstructionsMemory.m_mem[12]<=8'b00110100;
	InstructionsMemory.m_mem[13]<=8'b00100000;
	InstructionsMemory.m_mem[14]<=8'b00111011;
	InstructionsMemory.m_mem[15]<=8'b01010000;
	InstructionsMemory.m_mem[16]<=8'b00111100;
	InstructionsMemory.m_mem[17]<=8'b01100000;
	InstructionsMemory.m_mem[18]<=8'b11000111;
	InstructionsMemory.m_mem[19]<=8'b00010010;
	InstructionsMemory.m_mem[20]<=8'b11001000;
	InstructionsMemory.m_mem[21]<=8'b00010110;
	InstructionsMemory.m_mem[22]<=8'b11100111;
	InstructionsMemory.m_mem[23]<=8'b00000111;
	InstructionsMemory.m_mem[24]<=8'b11101000;
	InstructionsMemory.m_mem[25]<=8'b00001000;
	InstructionsMemory.m_mem[26]<=8'b11010010;
	InstructionsMemory.m_mem[27]<=8'b10001010;
	InstructionsMemory.m_mem[28]<=8'b10110010;
	InstructionsMemory.m_mem[29]<=8'b00000000;
	InstructionsMemory.m_mem[30]<=8'b00110100;
	InstructionsMemory.m_mem[31]<=8'b00100000;
	InstructionsMemory.m_mem[32]<=8'b00111011;
	InstructionsMemory.m_mem[33]<=8'b01011011;
	InstructionsMemory.m_mem[34]<=8'b00111100;
	InstructionsMemory.m_mem[35]<=8'b01101100;
	InstructionsMemory.m_mem[36]<=8'b11000111;
	InstructionsMemory.m_mem[37]<=8'b00010011;
	InstructionsMemory.m_mem[38]<=8'b11001000;
	InstructionsMemory.m_mem[39]<=8'b00010111;
	InstructionsMemory.m_mem[40]<=8'b11100111;
	InstructionsMemory.m_mem[41]<=8'b00000111;
	InstructionsMemory.m_mem[42]<=8'b11101000;
	InstructionsMemory.m_mem[43]<=8'b00001000;
	InstructionsMemory.m_mem[44]<=8'b11010010;
	InstructionsMemory.m_mem[45]<=8'b10001010;
	InstructionsMemory.m_mem[46]<=8'b10110010;
	InstructionsMemory.m_mem[47]<=8'b00000000;
	InstructionsMemory.m_mem[48]<=8'b00110100;
	InstructionsMemory.m_mem[49]<=8'b00100000;
	InstructionsMemory.m_mem[50]<=8'b00111011;
	InstructionsMemory.m_mem[51]<=8'b01011011;
	InstructionsMemory.m_mem[52]<=8'b00111100;
	InstructionsMemory.m_mem[53]<=8'b01101100;
	InstructionsMemory.m_mem[54]<=8'b11000111;
	InstructionsMemory.m_mem[55]<=8'b00010100;
	InstructionsMemory.m_mem[56]<=8'b11001000;
	InstructionsMemory.m_mem[57]<=8'b00011000;
	InstructionsMemory.m_mem[58]<=8'b11100111;
	InstructionsMemory.m_mem[59]<=8'b00000111;
	InstructionsMemory.m_mem[60]<=8'b11101000;
	InstructionsMemory.m_mem[61]<=8'b00001000;
	InstructionsMemory.m_mem[62]<=8'b11010010;
	InstructionsMemory.m_mem[63]<=8'b10001010;
	InstructionsMemory.m_mem[64]<=8'b10110010;
	InstructionsMemory.m_mem[65]<=8'b00000000;
	InstructionsMemory.m_mem[66]<=8'b00110100;
	InstructionsMemory.m_mem[67]<=8'b00100000;
	InstructionsMemory.m_mem[68]<=8'b00111100;
	InstructionsMemory.m_mem[69]<=8'b01101100;
	InstructionsMemory.m_mem[70]<=8'b00111011;
	InstructionsMemory.m_mem[71]<=8'b01011011;
	InstructionsMemory.m_mem[72]<=8'b11011101;
	InstructionsMemory.m_mem[73]<=8'b00000000;
	InstructionsMemory.m_mem[74]<=8'b11001110;
	InstructionsMemory.m_mem[75]<=8'b00000000;
	InstructionsMemory.m_mem[76]<=8'b11010010;
	InstructionsMemory.m_mem[77]<=8'b00001000;
	InstructionsMemory.m_mem[78]<=8'b10000010;
	InstructionsMemory.m_mem[79]<=8'b11010010;
	InstructionsMemory.m_mem[80]<=8'b11010010;
	InstructionsMemory.m_mem[81]<=8'b10000100;
	InstructionsMemory.m_mem[82]<=8'b00010010;
	InstructionsMemory.m_mem[83]<=8'b00000010;
	InstructionsMemory.m_mem[84]<=8'b11010010;
	InstructionsMemory.m_mem[85]<=8'b00000001;
	InstructionsMemory.m_mem[86]<=8'b01000011;
	InstructionsMemory.m_mem[87]<=8'b00110010;
	InstructionsMemory.m_mem[88]<=8'b11111101;
	InstructionsMemory.m_mem[89]<=8'b00000011;
	InstructionsMemory.m_mem[90]<=8'b11010010;
	InstructionsMemory.m_mem[91]<=8'b00000001;
	InstructionsMemory.m_mem[92]<=8'b01000011;
	InstructionsMemory.m_mem[93]<=8'b00110010;
	InstructionsMemory.m_mem[94]<=8'b11111110;
	InstructionsMemory.m_mem[95]<=8'b00000011;
	InstructionsMemory.m_mem[96]<=8'b11101101;
	InstructionsMemory.m_mem[97]<=8'b00001110;
	InstructionsMemory.m_mem[98]<=8'b11101110;
	InstructionsMemory.m_mem[99]<=8'b00011110;
	InstructionsMemory.m_mem[100]<=8'b01001101;
	InstructionsMemory.m_mem[101]<=8'b11001101;
	InstructionsMemory.m_mem[102]<=8'b01001110;
	InstructionsMemory.m_mem[103]<=8'b10111110;
	InstructionsMemory.m_mem[104]<=8'b00110010;
	InstructionsMemory.m_mem[105]<=8'b11011110;
	InstructionsMemory.m_mem[106]<=8'b11101110;
	InstructionsMemory.m_mem[107]<=8'b00000011;
	InstructionsMemory.m_mem[108]<=8'b11010010;
	InstructionsMemory.m_mem[109]<=8'b00000001;
	InstructionsMemory.m_mem[110]<=8'b00110011;
	InstructionsMemory.m_mem[111]<=8'b00110010;
	InstructionsMemory.m_mem[112]<=8'b11101101;
	InstructionsMemory.m_mem[113]<=8'b00000011;
	InstructionsMemory.m_mem[114]<=8'b11010010;
	InstructionsMemory.m_mem[115]<=8'b00000001;
	InstructionsMemory.m_mem[116]<=8'b00110011;
	InstructionsMemory.m_mem[117]<=8'b00110010;
	InstructionsMemory.m_mem[118]<=8'b11010010;
	InstructionsMemory.m_mem[119]<=8'b10000100;
	InstructionsMemory.m_mem[120]<=8'b00010000;
	InstructionsMemory.m_mem[121]<=8'b00100010;
	InstructionsMemory.m_mem[122]<=8'b11010010;
	InstructionsMemory.m_mem[123]<=8'b00000001;
	InstructionsMemory.m_mem[124]<=8'b00111101;
	InstructionsMemory.m_mem[125]<=8'b11010010;
	InstructionsMemory.m_mem[126]<=8'b11010010;
	InstructionsMemory.m_mem[127]<=8'b00000010;
	InstructionsMemory.m_mem[128]<=8'b00111110;
	InstructionsMemory.m_mem[129]<=8'b11100010;
	InstructionsMemory.m_mem[130]<=8'b10110000;
	InstructionsMemory.m_mem[131]<=8'b01001100;
	InstructionsMemory.m_mem[132]<=8'b11010010;
	InstructionsMemory.m_mem[133]<=8'b00000001;
	InstructionsMemory.m_mem[134]<=8'b00111101;
	InstructionsMemory.m_mem[135]<=8'b11010010;
	InstructionsMemory.m_mem[136]<=8'b00000001;
	InstructionsMemory.m_mem[137]<=8'b00000000;
	InstructionsMemory.m_mem[138]<=8'b11010010;
	InstructionsMemory.m_mem[139]<=8'b00000001;
	InstructionsMemory.m_mem[140]<=8'b01000011;
	InstructionsMemory.m_mem[141]<=8'b00110010;
	InstructionsMemory.m_mem[142]<=8'b11111011;
	InstructionsMemory.m_mem[143]<=8'b00000011;
	InstructionsMemory.m_mem[144]<=8'b11010010;
	InstructionsMemory.m_mem[145]<=8'b00000001;
	InstructionsMemory.m_mem[146]<=8'b01000011;
	InstructionsMemory.m_mem[147]<=8'b00110010;
	InstructionsMemory.m_mem[148]<=8'b11111100;
	InstructionsMemory.m_mem[149]<=8'b00000011;
	InstructionsMemory.m_mem[150]<=8'b10001011;
	InstructionsMemory.m_mem[151]<=8'b01111000;
	InstructionsMemory.m_mem[152]<=8'b11010010;
	InstructionsMemory.m_mem[153]<=8'b10100010;
	InstructionsMemory.m_mem[154]<=8'b00011011;
	InstructionsMemory.m_mem[155]<=8'b00000010;
	InstructionsMemory.m_mem[156]<=8'b00111011;
	InstructionsMemory.m_mem[157]<=8'b01110000;
	InstructionsMemory.m_mem[158]<=8'b00111100;
	InstructionsMemory.m_mem[159]<=8'b10000000;
	InstructionsMemory.m_mem[160]<=8'b10110000;
	InstructionsMemory.m_mem[161]<=8'b10100110;
	InstructionsMemory.m_mem[162]<=8'b00111011;
	InstructionsMemory.m_mem[163]<=8'b10000000;
	InstructionsMemory.m_mem[164]<=8'b00111100;
	InstructionsMemory.m_mem[165]<=8'b01110000;
	InstructionsMemory.m_mem[166]<=8'b11010101;
	InstructionsMemory.m_mem[167]<=8'b00000000;
	InstructionsMemory.m_mem[168]<=8'b11010110;
	InstructionsMemory.m_mem[169]<=8'b00000000;
	InstructionsMemory.m_mem[170]<=8'b11010010;
	InstructionsMemory.m_mem[171]<=8'b00000000;
	InstructionsMemory.m_mem[172]<=8'b10000010;
	InstructionsMemory.m_mem[173]<=8'b10110010;
	InstructionsMemory.m_mem[174]<=8'b01110010;
	InstructionsMemory.m_mem[175]<=8'b00100000;
	InstructionsMemory.m_mem[176]<=8'b11010010;
	InstructionsMemory.m_mem[177]<=8'b11000010;
	InstructionsMemory.m_mem[178]<=8'b00010010;
	InstructionsMemory.m_mem[179]<=8'b00000010;
	InstructionsMemory.m_mem[180]<=8'b00110101;
	InstructionsMemory.m_mem[181]<=8'b01011100;
	InstructionsMemory.m_mem[182]<=8'b11010111;
	InstructionsMemory.m_mem[183]<=8'b00000010;
	InstructionsMemory.m_mem[184]<=8'b11010010;
	InstructionsMemory.m_mem[185]<=8'b00000001;
	InstructionsMemory.m_mem[186]<=8'b00111011;
	InstructionsMemory.m_mem[187]<=8'b10110010;
	InstructionsMemory.m_mem[188]<=8'b11010010;
	InstructionsMemory.m_mem[189]<=8'b11010000;
	InstructionsMemory.m_mem[190]<=8'b00100001;
	InstructionsMemory.m_mem[191]<=8'b01110010;
	InstructionsMemory.m_mem[192]<=8'b10110000;
	InstructionsMemory.m_mem[193]<=8'b10101010;
	InstructionsMemory.m_mem[194]<=8'b11101100;
	InstructionsMemory.m_mem[195]<=8'b00000011;
	InstructionsMemory.m_mem[196]<=8'b11010010;
	InstructionsMemory.m_mem[197]<=8'b00000001;
	InstructionsMemory.m_mem[198]<=8'b00110011;
	InstructionsMemory.m_mem[199]<=8'b00110010;
	InstructionsMemory.m_mem[200]<=8'b11101011;
	InstructionsMemory.m_mem[201]<=8'b00000011;
	InstructionsMemory.m_mem[202]<=8'b11010010;
	InstructionsMemory.m_mem[203]<=8'b00000001;
	InstructionsMemory.m_mem[204]<=8'b00110011;
	InstructionsMemory.m_mem[205]<=8'b00110010;
	InstructionsMemory.m_mem[206]<=8'b10110100;
	InstructionsMemory.m_mem[207]<=8'b00000000;
	InstructionsMemory.m_mem[208]<=8'b11010010;
	InstructionsMemory.m_mem[209]<=8'b00000001;
	InstructionsMemory.m_mem[210]<=8'b00110110;
	InstructionsMemory.m_mem[211]<=8'b01100010;
	InstructionsMemory.m_mem[212]<=8'b10110000;
	InstructionsMemory.m_mem[213]<=8'b10101010;
	end
end
endmodule
